module main();

always @(posedge clock)
begin
  integer i;
  for(i=0; i<NUM_ROUTER; i=i+1)
  begin
    
  end
end

endmodule